module hashing();
endmodule